

module UART_Receiver (
    input wire clk,               // Clock input
    input wire rst,               // Reset input
    input wire rx,                // UART receive data
    output reg [7:0] data_out,    // 8-bit data outputs
    output reg crc_error          // CRC error flag
);

    localparam clks_per_bit = 1042; // Clock cycles per bit
    // State definitions for FSM
    localparam RX_IDLE       = 3'b000, // Receiver stay idle when rx = 1
               RX_START      = 3'b001, //  
               RX_DATA_TX    = 3'b010,  
               RX_CRC        = 3'b011,
               RX_STOP       = 3'b100;

    
    reg [2:0] rx_state = RX_IDLE;    // Current state of the FSM
    reg [2:0] bit_index;           // Bit index for data reception
    reg [12:0]clk_count;           // Clock count for baud rate
    reg [7:0] data_reg;            // Register to hold received data
    
    reg r_Rx_Data_R = 1'b1;
    reg r_data = 1'b1;
	 
    reg [3:0] crc_reg;             // Register to hold received 4-bit CRC code
    reg [3:0] computed_crc;        // Computed 4-bit CRC for verification
    reg [4:0] polynomial = 5'b10011;           // Polynomial x^4 + x + 1 (binary: 10011)
	 
	 // Compute CRC on positive edge of `tx_start`
    always @(posedge clk) begin
	 
        if (rx_state == RX_STOP) begin
           computed_crc <= CHECK_CRC({data_reg,crc_reg});
        end
		
    end
   
	 // Task to check for error 
	 function [3:0] CHECK_CRC;
        input [11:0] data_crc;  // 12-bit input: 8-bit data + 4-bit CRC
        reg [3:0] remainder;
        begin
            // Step-by-step manual XOR operations to simulate polynomial division
            remainder[3] = data_crc[11] ^ data_crc[7] ^ data_crc[4] ^ data_crc[3] ^ data_crc[0];
            remainder[2] = data_crc[10] ^ data_crc[6] ^ data_crc[3];
            remainder[1] = data_crc[9] ^ data_crc[5] ^ data_crc[2];
            remainder[0] = data_crc[8] ^ data_crc[4] ^ data_crc[1] ^ data_crc[0];

            // Check if remainder is zero
            CHECK_CRC = remainder;
				
        end
    endfunction
	 
    // Purpose: Double-register the incoming data.
    always @(posedge clk) begin
        r_Rx_Data_R <= rx;
        r_data <= r_Rx_Data_R;
		  end
    
    always @(posedge clk) begin
	 
        if (rst) begin
            rx_state <= RX_IDLE;
            clk_count <= 0;
            bit_index <= 0;
            crc_error <= 0;
				data_out <= 8'b0;
        end 
		  
		  else begin  
				case (rx_state)
                RX_IDLE: begin
                    crc_error <= 0;
                    clk_count <= 0;
                    bit_index <= 0;
						  
                    if (r_data == 1'b0) begin
                        rx_state <= RX_START;
						  end
						  end // END CASE: FOR RX_IDLE
                 
					 RX_START : begin
							if(clk_count < (clks_per_bit)/2) begin
							   clk_count <= clk_count + 1;
								end
								else begin
								if (r_data == 1'b0)begin
									bit_index <= 0;
									clk_count <= 0;
									rx_state <= RX_DATA_TX;
									end
									end
									end // END CASE FOR RX_START
									
					 
					 RX_DATA_TX : begin
						if (clk_count < clks_per_bit) begin
							 clk_count<= clk_count + 1;

							end
						
						else begin
								 
										data_reg[bit_index] <= r_data;
                 
									 // Check if we have received all bits
										if (bit_index < 7)
										begin
										  clk_count <= 0;
										  bit_index <= bit_index + 1;
										 rx_state   <=  RX_DATA_TX;
										end
										
									 else
										begin
										  clk_count <=0;
										  bit_index <= 0;
										  rx_state   <= RX_CRC;
										end
								  end
							 end // case: RX_DATA_TX
			 
			       RX_CRC : begin
			       
					 if (clk_count < clks_per_bit) begin
							 clk_count <= clk_count + 1;
							end
							
							else begin 
								 crc_reg[bit_index] <= r_data;
                                                      
							 // Check if we have received all bits
								if (bit_index < 3)
								begin
								  clk_count <= 0;
								  bit_index <= bit_index + 1;
								  rx_state   <=  RX_CRC;
								end
								
							 else
								begin
								  bit_index <= 0;
								  clk_count <= 0;
								  rx_state   <= RX_STOP;
								end
						  end
					 end // case: RX_CRC 
					 
																
				RX_STOP : begin
				     // Compute CRC

                 // Wait clks_per_bit clock cycles for Stop bit to finish
						if (clk_count < clks_per_bit)
							begin
								clk_count <= clk_count + 1;
								rx_state <= RX_STOP;
							end
					
					  	 else
							begin
							  
								if(r_data == 1'b1) begin  // Stop bit check
									if(computed_crc == 4'b0000) begin
										crc_error <= 1'b0;  // CRC mismatch error
										data_out <= data_reg;
										rx_state <= RX_IDLE;
										end
										
									else begin
										crc_error <= 1'b1; // No error
										data_out <= 8'b00000000;
										rx_state <= RX_IDLE;
										end
										end
			          	 end 
			             end // case:RX_STOP
							 
							default: 
								rx_state <= RX_IDLE;
						   endcase
					end // END OF CASE STATEMENT
				end // END OF ALWAYS 	
				
endmodule 

